-- Ifetch module (provides the PC and instruction 
--memory for the MIPS computer)
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
LIBRARY altera_mf;
USE altera_mf.altera_mf_components.all;

ENTITY Ifetch IS
	PORT(	SIGNAL Instruction 		: OUT	STD_LOGIC_VECTOR( 31 DOWNTO 0 );
        	SIGNAL PC_plus_4_out 	: OUT	STD_LOGIC_VECTOR( 9 DOWNTO 0 );
        	SIGNAL Add_result 		: IN 	STD_LOGIC_VECTOR( 7 DOWNTO 0 );
        	SIGNAL BranchEQ 		: IN 	STD_LOGIC;
        	SIGNAL BranchNEQ 		: IN 	STD_LOGIC;
        	SIGNAL Zero,j,jr 			: IN 	STD_LOGIC;
      		SIGNAL PC_out 			: OUT	STD_LOGIC_VECTOR( 9 DOWNTO 0 );
        	SIGNAL clock, reset 	: IN 	STD_LOGIC;
			SIGNAL ALU_result_jr 		: IN 	STD_LOGIC_VECTOR( 7 DOWNTO 0 ));
END Ifetch;

ARCHITECTURE behavior OF Ifetch IS
	SIGNAL PC, PC_plus_4, Mem_Addr : STD_LOGIC_VECTOR( 9 DOWNTO 0 );
	SIGNAL next_PC,jumpaddress : STD_LOGIC_VECTOR( 7 DOWNTO 0 );
	SIGNAL Instruction_sig 		: 	STD_LOGIC_VECTOR( 31 DOWNTO 0 );
BEGIN
						--ROM for Instruction Memory
inst_memory: altsyncram
	
	GENERIC MAP (
		operation_mode => "ROM",
		width_a => 32,
		widthad_a => 10,
		lpm_type => "altsyncram",
		outdata_reg_a => "UNREGISTERED",
		init_file => "C:\Users\TalKa\Documents\GitHub\Task3newest\MIPS Quartus\text.hex",
		intended_device_family => "Cyclone"
	)
	PORT MAP (
		clock0      => clock,
		address_a 	=> Mem_Addr, 
		q_a 		=> Instruction_sig );
		
		Instruction <= Instruction_sig;
		jumpaddress(7 downto 0)<= Instruction_sig( 7 DOWNTO 0);
		
					-- Instructions always start on word address - not byte
		PC(1 DOWNTO 0) <= "00";
					-- copy output signals - allows read inside module
		PC_out 			<= PC;
		PC_plus_4_out 	<= PC_plus_4;
						-- send address to inst. memory address register
						
		Mem_Addr <=    Next_PC & "00" ; --Quartos				
		-- Mem_Addr <=  "00" & Next_PC    ; --MODELSIM

						-- Adder to increment PC by 4        
      	PC_plus_4( 9 DOWNTO 2 )  <= PC( 9 DOWNTO 2 ) + 1;
       	PC_plus_4( 1 DOWNTO 0 )  <= "00";
						-- Mux to select Branch Address or PC + 4        
		Next_PC  <= X"00" WHEN Reset = '1' ELSE -- for reset
			ALU_result_jr  WHEN jr = '1' ELSE -- for Jr
			Add_result  WHEN ( ( BranchEQ = '1' ) AND ( Zero = '1' ) ) ELSE -- for BEQ
			Add_result  WHEN ( ( BranchNEQ = '1' ) AND ( Zero = '0' ) ) ELSE -- for BNE
			jumpaddress	WHEN (j ='1') ELSE -- for jump
			PC_plus_4( 9 DOWNTO 2 ); -- normal state, pc + 4
	PROCESS
		BEGIN
			WAIT UNTIL ( clock'EVENT ) AND ( clock = '1' );
			IF reset = '1' THEN
				   PC( 9 DOWNTO 2) <= "00000000" ; 
			ELSE 
				   PC( 9 DOWNTO 2 ) <= next_PC;
			END IF;
	END PROCESS;
END behavior;


